module alchitry_tb_top;

endmodule : alchitry_tb_top
