module alchitry_top;


endmodule : alchitry_top
